mailbox gen2bfm=new();
mailbox mon2cov=new();
mailbox mon2sbd=new();
parameter n=3;
static int num_matches;  // If a varaiable gets static then it can be accessed everywhere.
static int num_miss_matches;
static int  count=3;
