`include "common.sv"
`include "interface.sv"
`include "transaction.sv"
`include "binary2grey_gen.sv"
`include "binary2grey_bfm.sv"
`include "binary2grey_mon.sv"
`include "binary2grey_cov.sv"
`include "binary2grey_agent.sv"
`include "binary2grey_sbd.sv"
`include "binary2grey_env.sv"
`include "module_top.sv"
