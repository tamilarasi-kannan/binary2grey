interface binary2grey_int();
  bit [n-1:0]binary,grey;
endinterface
